----------------------------------------------------------------------------------------------------
-- Engineer: T�th �d�m Raymond
-- Advisor: Dr. Horv�th P�ter

-- University: Budapesti M�szaki �s Gazdas�gtudom�nyi Egyetem
-- Faculty: Villamosm�rn�ki �s Informatikai Kar
-- Department: Elektronikus Eszk�z�k Tansz�k

-- Semester: 2019/20/2

-- Design Name: �jrafelhaszn�lhat� mem�riamodul nagymegb�zhat�s�g� rendszerekhez
-- Module Name:

-- Description: 

----------------------------------------------------------------------------------------------------


library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.math_real.all;


entity counter is
    generic(
        -- clock: 100 MHz
        
        -- prescaler counts to seconds (depends on the clock)
        -- prescaler: 2**size
        prescaler_size: integer := 17;
        
        -- timer counts to hours (depends on the user)
        --timer: 2**size
        timer_size: integer := 9
    );
    port(
        clk: in std_logic;
        rst_n: in std_logic;
        input_idle: in std_logic;
        force: in std_logic;
        wakeup: out std_logic
    );
end counter;

architecture rtl of counter is

    signal prescaler: std_logic_vector((prescaler_size-1) downto 0) := (others => '1');
    signal timer: std_logic_vector((timer_size-1) downto 0) := (others => '1');

begin

    L_TIMER: process(clk,rst_n)
    begin
        if(rst_n = '0') then
            prescaler <= (others => '1');
            timer <= (others => '1');
        elsif(rising_edge(clk)) then
            if(force = '1') then
                prescaler <= (others => '1');
                timer <= (others => '1');
            elsif(input_idle = '1') then
                prescaler <= std_logic_vector(unsigned(prescaler) - 1);
                if(unsigned(prescaler) = 0) then
                    timer <= std_logic_vector(unsigned(timer) - 1);
                end if;
            end if;
        end if;
    end process;
    wakeup <= '1' when ((unsigned(prescaler) = 0) and (unsigned(timer) = 0));

end rtl;
